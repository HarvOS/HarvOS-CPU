// bus_if.sv (minimal) — Interfaces moved to standalone files.
// harvos_imem_if is defined in harvos_imem_if.sv
// harvos_dmem_if is defined in harvos_dmem_if.sv
// This file intentionally left minimal to avoid redefinitions during synthesis.
